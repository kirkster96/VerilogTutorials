module and2_v(y,b,a);
	output y;       // module output
	input  b,a;     // module input
	assign y = a&b; // continuous assignment
endmodule
