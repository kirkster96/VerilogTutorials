// (C) 2001-2017 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// seq.v

// This file was auto-generated from qsys_sequencer_110_hw.tcl.  If you edit it your changes
// will probably be lost.
// 
// Generated using ACDS version 11.1 147 at 2011.09.14.12:07:16

`timescale 1 ps / 1 ps
module seq (
		input  wire        avl_clk,                 //          avl_clk.clk
		input  wire        avl_reset_n,             //        avl_reset.reset_n
		input  wire        apb_clk,                 //          apb_clk.clk
		input  wire        apb_reset_n,             //        apb_reset.reset_n
		output wire [31:0] prdata,                  //        apb_slave.prdata
		output wire        pready,                  //                 .pready
		output wire        pslverr,                 //                 .pslverr
		input  wire [31:0] pwdata,                  //                 .pwdata
		input  wire        pwrite,                  //                 .pwrite
		input  wire        penable,                 //                 .penable
		input  wire        psel,                    //                 .psel
		input  wire [31:0] paddr,                   //                 .paddr
		input  wire        mmr_avl_waitrequest,     //          mmr_avl.waitrequest
		input  wire [31:0] mmr_avl_readdata,        //                 .readdata
		input  wire        mmr_avl_readdatavalid,   //                 .readdatavalid
		output wire        mmr_avl_burstcount,      //                 .burstcount
		output wire [31:0] mmr_avl_writedata,       //                 .writedata
		output wire [7:0]  mmr_avl_address,         //                 .address
		output wire        mmr_avl_write,           //                 .write
		output wire        mmr_avl_read,            //                 .read
//		output wire [3:0]  mmr_avl_be,              //                 .byteenable
		output wire        mmr_avl_debugaccess,     //                 .debugaccess
		output wire [15:0] avl_address,             //              avl.address
		output wire        avl_read,                //                 .read
		input  wire [31:0] avl_readdata,            //                 .readdata
		output wire        avl_write,               //                 .write
		output wire [31:0] avl_writedata,           //                 .writedata
		input  wire        avl_waitrequest,         //                 .waitrequest
		output wire        scc_data,                //              scc.scc_data
		output wire [4:0]  scc_dqs_ena,             //                 .scc_dqs_ena
		output wire [4:0]  scc_dqsb_ena,             //                 .scc_dqs_ena
		output wire [4:0]  scc_dqs_io_ena,          //                 .scc_dqs_io_ena
		output wire [39:0] scc_dq_ena,              //                 .scc_dq_ena
		output wire [4:0]  scc_dm_ena,              //                 .scc_dm_ena
		output wire        scc_upd,                 //                 .scc_upd
		input  wire [4:0]  capture_strobe_tracking, //                 .capture_strobe_tracking
		input  wire        afi_init_req,            // afi_init_cal_req.afi_init_req
		input  wire        afi_cal_req,             //                 .afi_cal_req
//		input  wire        scc_clk,                 //          scc_clk.clk
		output wire [4:0]  scc_clk_out,
//		input  wire        reset_n_scc_clk,         //        scc_reset.reset_n
		output wire [1:0]  afi_seq_busy,            //          trk_afi.afi_seq_busy
		input  wire [1:0]  afi_ctl_long_idle,       //                 .afi_ctl_long_idle
		input  wire [1:0]  afi_ctl_refresh_done,    //                 .afi_ctl_refresh_done
		
		//debug signals
		output wire [58:0] debug_hphy_reg,
		output wire [42:0] debug_hphy_comb

		
	);
	
	//debug signals
	wire [18:0] debug_hphy_reg_scc;
	wire [12:0] debug_hphy_comb_scc;

	wire [ 2:0] debug_hphy_reg_reg;
	wire        debug_hphy_comb_reg;

	wire [24:0] debug_hphy_reg_trck;
	wire [ 1:0] debug_hphy_comb_trck;

	wire [ 8:0] debug_hphy_reg_apb2avl;
	wire        debug_hphy_comb_apb2avl;

	wire [18:0] debug_hphy_comb_decompress;

	wire  [2:0] debug_hphy_reg_clk_crossing;
	wire  [6:0] debug_hphy_comb_clk_crossing;
 

	wire         apb2avalon_bridge_inst_avalon_master_waitrequest;                                                 // apb2avalon_bridge_inst_avalon_master_translator:av_waitrequest -> apb2avalon_bridge_inst:av_waitrequest
	wire  [31:0] apb2avalon_bridge_inst_avalon_master_writedata;                                                   // apb2avalon_bridge_inst:av_writedata -> apb2avalon_bridge_inst_avalon_master_translator:av_writedata
	wire  [31:0] apb2avalon_bridge_inst_avalon_master_address;                                                     // apb2avalon_bridge_inst:av_addr -> apb2avalon_bridge_inst_avalon_master_translator:av_address
	wire         apb2avalon_bridge_inst_avalon_master_write;                                                       // apb2avalon_bridge_inst:av_write -> apb2avalon_bridge_inst_avalon_master_translator:av_write
	wire         apb2avalon_bridge_inst_avalon_master_read;                                                        // apb2avalon_bridge_inst:av_read -> apb2avalon_bridge_inst_avalon_master_translator:av_read
	wire  [31:0] apb2avalon_bridge_inst_avalon_master_readdata;                                                    // apb2avalon_bridge_inst_avalon_master_translator:av_readdata -> apb2avalon_bridge_inst:av_readdata
	wire   [3:0] apb2avalon_bridge_inst_avalon_master_byteenable;                                                  // apb2avalon_bridge_inst:av_byteenable -> apb2avalon_bridge_inst_avalon_master_translator:av_byteenable
	wire         apb2avalon_bridge_inst_avalon_master_readdatavalid;                                               // apb2avalon_bridge_inst_avalon_master_translator:av_readdatavalid -> apb2avalon_bridge_inst:av_rdata_valid
	wire         apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_waitrequest;            // seq_hhp_decompress_bridge_s0_translator:uav_waitrequest -> apb2avalon_bridge_inst_avalon_master_translator:uav_waitrequest
	wire   [2:0] apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_burstcount;             // apb2avalon_bridge_inst_avalon_master_translator:uav_burstcount -> seq_hhp_decompress_bridge_s0_translator:uav_burstcount
	wire  [31:0] apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_writedata;              // apb2avalon_bridge_inst_avalon_master_translator:uav_writedata -> seq_hhp_decompress_bridge_s0_translator:uav_writedata
	wire  [31:0] apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_address;                // apb2avalon_bridge_inst_avalon_master_translator:uav_address -> seq_hhp_decompress_bridge_s0_translator:uav_address
	wire         apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_lock;                   // apb2avalon_bridge_inst_avalon_master_translator:uav_lock -> seq_hhp_decompress_bridge_s0_translator:uav_lock
	wire         apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_write;                  // apb2avalon_bridge_inst_avalon_master_translator:uav_write -> seq_hhp_decompress_bridge_s0_translator:uav_write
	wire         apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_read;                   // apb2avalon_bridge_inst_avalon_master_translator:uav_read -> seq_hhp_decompress_bridge_s0_translator:uav_read
	wire  [31:0] apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_readdata;               // seq_hhp_decompress_bridge_s0_translator:uav_readdata -> apb2avalon_bridge_inst_avalon_master_translator:uav_readdata
	wire         apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_debugaccess;            // apb2avalon_bridge_inst_avalon_master_translator:uav_debugaccess -> seq_hhp_decompress_bridge_s0_translator:uav_debugaccess
	wire   [3:0] apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_byteenable;             // apb2avalon_bridge_inst_avalon_master_translator:uav_byteenable -> seq_hhp_decompress_bridge_s0_translator:uav_byteenable
	wire         apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_readdatavalid;          // seq_hhp_decompress_bridge_s0_translator:uav_readdatavalid -> apb2avalon_bridge_inst_avalon_master_translator:uav_readdatavalid
	wire         seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                              // seq_hhp_decompress_bridge:s0_waitrequest -> seq_hhp_decompress_bridge_s0_translator:av_waitrequest
	wire  [31:0] seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_writedata;                                // seq_hhp_decompress_bridge_s0_translator:av_writedata -> seq_hhp_decompress_bridge:s0_writedata
	wire  [31:0] seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_address;                                  // seq_hhp_decompress_bridge_s0_translator:av_address -> seq_hhp_decompress_bridge:s0_address
	wire         seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_write;                                    // seq_hhp_decompress_bridge_s0_translator:av_write -> seq_hhp_decompress_bridge:s0_write
	wire         seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_read;                                     // seq_hhp_decompress_bridge_s0_translator:av_read -> seq_hhp_decompress_bridge:s0_read
	wire  [31:0] seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_readdata;                                 // seq_hhp_decompress_bridge:s0_readdata -> seq_hhp_decompress_bridge_s0_translator:av_readdata
	wire         seq_hhp_decompress_bridge_m0_waitrequest;                                                             // seq_hhp_decompress_bridge_m0_translator:av_waitrequest -> seq_hhp_decompress_bridge:m0_waitrequest
	wire  [31:0] seq_hhp_decompress_bridge_m0_writedata;                                                               // seq_hhp_decompress_bridge:m0_writedata -> seq_hhp_decompress_bridge_m0_translator:av_writedata
	wire  [31:0] seq_hhp_decompress_bridge_m0_address;                                                                 // seq_hhp_decompress_bridge:m0_address -> seq_hhp_decompress_bridge_m0_translator:av_address
	wire         seq_hhp_decompress_bridge_m0_write;                                                                   // seq_hhp_decompress_bridge:m0_write -> seq_hhp_decompress_bridge_m0_translator:av_write
	wire         seq_hhp_decompress_bridge_m0_read;                                                                    // seq_hhp_decompress_bridge:m0_read -> seq_hhp_decompress_bridge_m0_translator:av_read
	wire  [31:0] seq_hhp_decompress_bridge_m0_readdata;                                                                // seq_hhp_decompress_bridge_m0_translator:av_readdata -> seq_hhp_decompress_bridge:m0_readdata
	wire         seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_waitrequest;                        // cpu_inst_s0_translator:uav_waitrequest -> seq_hhp_decompress_bridge_m0_translator:uav_waitrequest
	wire   [2:0] seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_burstcount;                         // seq_hhp_decompress_bridge_m0_translator:uav_burstcount -> cpu_inst_s0_translator:uav_burstcount
	wire  [31:0] seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_writedata;                          // seq_hhp_decompress_bridge_m0_translator:uav_writedata -> cpu_inst_s0_translator:uav_writedata
	wire  [31:0] seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_address;                            // seq_hhp_decompress_bridge_m0_translator:uav_address -> cpu_inst_s0_translator:uav_address
	wire         seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_lock;                               // seq_hhp_decompress_bridge_m0_translator:uav_lock -> cpu_inst_s0_translator:uav_lock
	wire         seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_write;                              // seq_hhp_decompress_bridge_m0_translator:uav_write -> cpu_inst_s0_translator:uav_write
	wire         seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_read;                               // seq_hhp_decompress_bridge_m0_translator:uav_read -> cpu_inst_s0_translator:uav_read
	wire  [31:0] seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_readdata;                           // cpu_inst_s0_translator:uav_readdata -> seq_hhp_decompress_bridge_m0_translator:uav_readdata
	wire         seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_debugaccess;                        // seq_hhp_decompress_bridge_m0_translator:uav_debugaccess -> cpu_inst_s0_translator:uav_debugaccess
	wire   [3:0] seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_byteenable;                         // seq_hhp_decompress_bridge_m0_translator:uav_byteenable -> cpu_inst_s0_translator:uav_byteenable
	wire         seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                      // cpu_inst_s0_translator:uav_readdatavalid -> seq_hhp_decompress_bridge_m0_translator:uav_readdatavalid
	wire         cpu_inst_s0_translator_avalon_anti_slave_0_waitrequest;                                           // cpu_inst:s0_waitrequest -> cpu_inst_s0_translator:av_waitrequest
	wire         cpu_inst_s0_translator_avalon_anti_slave_0_burstcount;                                            // cpu_inst_s0_translator:av_burstcount -> cpu_inst:s0_burstcount
	wire  [31:0] cpu_inst_s0_translator_avalon_anti_slave_0_writedata;                                             // cpu_inst_s0_translator:av_writedata -> cpu_inst:s0_writedata
	wire  [19:0] cpu_inst_s0_translator_avalon_anti_slave_0_address;                                               // cpu_inst_s0_translator:av_address -> cpu_inst:s0_address
	wire         cpu_inst_s0_translator_avalon_anti_slave_0_write;                                                 // cpu_inst_s0_translator:av_write -> cpu_inst:s0_write
	wire         cpu_inst_s0_translator_avalon_anti_slave_0_read;                                                  // cpu_inst_s0_translator:av_read -> cpu_inst:s0_read
	wire  [31:0] cpu_inst_s0_translator_avalon_anti_slave_0_readdata;                                              // cpu_inst:s0_readdata -> cpu_inst_s0_translator:av_readdata
	wire         cpu_inst_s0_translator_avalon_anti_slave_0_debugaccess;                                           // cpu_inst_s0_translator:av_debugaccess -> cpu_inst:s0_debugaccess
	wire         cpu_inst_s0_translator_avalon_anti_slave_0_readdatavalid;                                         // cpu_inst:s0_readdatavalid -> cpu_inst_s0_translator:av_readdatavalid
	wire   [3:0] cpu_inst_s0_translator_avalon_anti_slave_0_byteenable;                                            // cpu_inst_s0_translator:av_byteenable -> cpu_inst:s0_byteenable
	wire   [0:0] cpu_inst_m0_burstcount;                                                                           // cpu_inst:m0_burstcount -> cpu_inst_m0_translator:av_burstcount
	wire         cpu_inst_m0_waitrequest;                                                                          // cpu_inst_m0_translator:av_waitrequest -> cpu_inst:m0_waitrequest
	wire  [19:0] cpu_inst_m0_address;                                                                              // cpu_inst:m0_address -> cpu_inst_m0_translator:av_address
	wire  [31:0] cpu_inst_m0_writedata;                                                                            // cpu_inst:m0_writedata -> cpu_inst_m0_translator:av_writedata
	wire         cpu_inst_m0_write;                                                                                // cpu_inst:m0_write -> cpu_inst_m0_translator:av_write
	wire         cpu_inst_m0_read;                                                                                 // cpu_inst:m0_read -> cpu_inst_m0_translator:av_read
	wire  [31:0] cpu_inst_m0_readdata;                                                                             // cpu_inst_m0_translator:av_readdata -> cpu_inst:m0_readdata
	wire         cpu_inst_m0_debugaccess;                                                                          // cpu_inst:m0_debugaccess -> cpu_inst_m0_translator:av_debugaccess
	wire   [3:0] cpu_inst_m0_byteenable;                                                                           // cpu_inst:m0_byteenable -> cpu_inst_m0_translator:av_byteenable
	wire         cpu_inst_m0_readdatavalid;                                                                        // cpu_inst_m0_translator:av_readdatavalid -> cpu_inst:m0_readdatavalid
	wire         seq_trk_mgr_inst_avl_waitrequest;                                                           // seq_trk_mgr_inst_avl_translator:av_waitrequest -> seq_trk_mgr_inst:avl_waitrequest
	wire  [31:0] seq_trk_mgr_inst_avl_writedata;                                                             // seq_trk_mgr_inst:avl_writedata -> seq_trk_mgr_inst_avl_translator:av_writedata
	wire  [19:0] seq_trk_mgr_inst_avl_address;                                                               // seq_trk_mgr_inst:avl_address -> seq_trk_mgr_inst_avl_translator:av_address
	wire         seq_trk_mgr_inst_avl_write;                                                                 // seq_trk_mgr_inst:avl_write -> seq_trk_mgr_inst_avl_translator:av_write
	wire         seq_trk_mgr_inst_avl_read;                                                                  // seq_trk_mgr_inst:avl_read -> seq_trk_mgr_inst_avl_translator:av_read
	wire  [31:0] seq_trk_mgr_inst_avl_readdata;                                                              // seq_trk_mgr_inst_avl_translator:av_readdata -> seq_trk_mgr_inst:avl_readdata
	wire         mmr_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                         // mmr_bridge:s0_waitrequest -> mmr_bridge_s0_translator:av_waitrequest
	wire         mmr_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                          // mmr_bridge_s0_translator:av_burstcount -> mmr_bridge:s0_burstcount
	wire  [31:0] mmr_bridge_s0_translator_avalon_anti_slave_0_writedata;                                           // mmr_bridge_s0_translator:av_writedata -> mmr_bridge:s0_writedata
	wire   [7:0] mmr_bridge_s0_translator_avalon_anti_slave_0_address;                                             // mmr_bridge_s0_translator:av_address -> mmr_bridge:s0_address
	wire         mmr_bridge_s0_translator_avalon_anti_slave_0_write;                                               // mmr_bridge_s0_translator:av_write -> mmr_bridge:s0_write
	wire         mmr_bridge_s0_translator_avalon_anti_slave_0_read;                                                // mmr_bridge_s0_translator:av_read -> mmr_bridge:s0_read
	wire  [31:0] mmr_bridge_s0_translator_avalon_anti_slave_0_readdata;                                            // mmr_bridge:s0_readdata -> mmr_bridge_s0_translator:av_readdata
	wire         mmr_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                         // mmr_bridge_s0_translator:av_debugaccess -> mmr_bridge:s0_debugaccess
	wire         mmr_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                       // mmr_bridge:s0_readdatavalid -> mmr_bridge_s0_translator:av_readdatavalid
	wire   [3:0] mmr_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                          // mmr_bridge_s0_translator:av_byteenable -> mmr_bridge:s0_byteenable
	wire         hphy_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                        // hphy_bridge:s0_waitrequest -> hphy_bridge_s0_translator:av_waitrequest
	wire  [31:0] hphy_bridge_s0_translator_avalon_anti_slave_0_writedata;                                          // hphy_bridge_s0_translator:av_writedata -> hphy_bridge:s0_writedata
	wire  [15:0] hphy_bridge_s0_translator_avalon_anti_slave_0_address;                                            // hphy_bridge_s0_translator:av_address -> hphy_bridge:s0_address
	wire         hphy_bridge_s0_translator_avalon_anti_slave_0_write;                                              // hphy_bridge_s0_translator:av_write -> hphy_bridge:s0_write
	wire         hphy_bridge_s0_translator_avalon_anti_slave_0_read;                                               // hphy_bridge_s0_translator:av_read -> hphy_bridge:s0_read
	wire  [31:0] hphy_bridge_s0_translator_avalon_anti_slave_0_readdata;                                           // hphy_bridge:s0_readdata -> hphy_bridge_s0_translator:av_readdata
	wire         seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_waitrequest;                            // seq_scc_mgr_inst:avl_waitrequest -> seq_scc_mgr_inst_avl_translator:av_waitrequest
	wire  [31:0] seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_writedata;                              // seq_scc_mgr_inst_avl_translator:av_writedata -> seq_scc_mgr_inst:avl_writedata
	wire  [12:0] seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_address;                                // seq_scc_mgr_inst_avl_translator:av_address -> seq_scc_mgr_inst:avl_address
	wire         seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_write;                                  // seq_scc_mgr_inst_avl_translator:av_write -> seq_scc_mgr_inst:avl_write
	wire         seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_read;                                   // seq_scc_mgr_inst_avl_translator:av_read -> seq_scc_mgr_inst:avl_read
	wire  [31:0] seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_readdata;                               // seq_scc_mgr_inst:avl_readdata -> seq_scc_mgr_inst_avl_translator:av_readdata
	wire         seq_reg_file_inst_avl_translator_avalon_anti_slave_0_waitrequest;                           // seq_reg_file_inst:avl_waitrequest -> seq_reg_file_inst_avl_translator:av_waitrequest
	wire  [31:0] seq_reg_file_inst_avl_translator_avalon_anti_slave_0_writedata;                             // seq_reg_file_inst_avl_translator:av_writedata -> seq_reg_file_inst:avl_writedata
	wire  [12:0] seq_reg_file_inst_avl_translator_avalon_anti_slave_0_address;                               // seq_reg_file_inst_avl_translator:av_address -> seq_reg_file_inst:avl_address
	wire         seq_reg_file_inst_avl_translator_avalon_anti_slave_0_write;                                 // seq_reg_file_inst_avl_translator:av_write -> seq_reg_file_inst:avl_write
	wire         seq_reg_file_inst_avl_translator_avalon_anti_slave_0_read;                                  // seq_reg_file_inst_avl_translator:av_read -> seq_reg_file_inst:avl_read
	wire  [31:0] seq_reg_file_inst_avl_translator_avalon_anti_slave_0_readdata;                              // seq_reg_file_inst:avl_readdata -> seq_reg_file_inst_avl_translator:av_readdata
	wire   [3:0] seq_reg_file_inst_avl_translator_avalon_anti_slave_0_byteenable;                            // seq_reg_file_inst_avl_translator:av_byteenable -> seq_reg_file_inst:avl_be
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // seq_reg_file_inst_avl_translator:uav_waitrequest -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:m0_burstcount -> seq_reg_file_inst_avl_translator:uav_burstcount
	wire  [31:0] seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_writedata;               // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:m0_writedata -> seq_reg_file_inst_avl_translator:uav_writedata
	wire  [19:0] seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_address;                 // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:m0_address -> seq_reg_file_inst_avl_translator:uav_address
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_write;                   // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:m0_write -> seq_reg_file_inst_avl_translator:uav_write
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_lock;                    // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:m0_lock -> seq_reg_file_inst_avl_translator:uav_lock
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_read;                    // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:m0_read -> seq_reg_file_inst_avl_translator:uav_read
	wire  [31:0] seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdata;                // seq_reg_file_inst_avl_translator:uav_readdata -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // seq_reg_file_inst_avl_translator:uav_readdatavalid -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> seq_reg_file_inst_avl_translator:uav_debugaccess
	wire   [3:0] seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:m0_byteenable -> seq_reg_file_inst_avl_translator:uav_byteenable
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rf_source_valid -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [73:0] seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_data;             // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rf_source_data -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [73:0] seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_inst_m0_translator_avalon_universal_master_0_waitrequest;                                     // cpu_inst_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_inst_m0_translator:uav_waitrequest
	wire   [2:0] cpu_inst_m0_translator_avalon_universal_master_0_burstcount;                                      // cpu_inst_m0_translator:uav_burstcount -> cpu_inst_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_inst_m0_translator_avalon_universal_master_0_writedata;                                       // cpu_inst_m0_translator:uav_writedata -> cpu_inst_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire  [19:0] cpu_inst_m0_translator_avalon_universal_master_0_address;                                         // cpu_inst_m0_translator:uav_address -> cpu_inst_m0_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_inst_m0_translator_avalon_universal_master_0_lock;                                            // cpu_inst_m0_translator:uav_lock -> cpu_inst_m0_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_inst_m0_translator_avalon_universal_master_0_write;                                           // cpu_inst_m0_translator:uav_write -> cpu_inst_m0_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_inst_m0_translator_avalon_universal_master_0_read;                                            // cpu_inst_m0_translator:uav_read -> cpu_inst_m0_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_inst_m0_translator_avalon_universal_master_0_readdata;                                        // cpu_inst_m0_translator_avalon_universal_master_0_agent:av_readdata -> cpu_inst_m0_translator:uav_readdata
	wire         cpu_inst_m0_translator_avalon_universal_master_0_debugaccess;                                     // cpu_inst_m0_translator:uav_debugaccess -> cpu_inst_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_inst_m0_translator_avalon_universal_master_0_byteenable;                                      // cpu_inst_m0_translator:uav_byteenable -> cpu_inst_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_inst_m0_translator_avalon_universal_master_0_readdatavalid;                                   // cpu_inst_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_inst_m0_translator:uav_readdatavalid
	wire         seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_waitrequest;                      // seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:av_waitrequest -> seq_trk_mgr_inst_avl_translator:uav_waitrequest
	wire   [2:0] seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_burstcount;                       // seq_trk_mgr_inst_avl_translator:uav_burstcount -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_writedata;                        // seq_trk_mgr_inst_avl_translator:uav_writedata -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:av_writedata
	wire  [19:0] seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_address;                          // seq_trk_mgr_inst_avl_translator:uav_address -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:av_address
	wire         seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_lock;                             // seq_trk_mgr_inst_avl_translator:uav_lock -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:av_lock
	wire         seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_write;                            // seq_trk_mgr_inst_avl_translator:uav_write -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:av_write
	wire         seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_read;                             // seq_trk_mgr_inst_avl_translator:uav_read -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_readdata;                         // seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:av_readdata -> seq_trk_mgr_inst_avl_translator:uav_readdata
	wire         seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_debugaccess;                      // seq_trk_mgr_inst_avl_translator:uav_debugaccess -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_byteenable;                       // seq_trk_mgr_inst_avl_translator:uav_byteenable -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:av_byteenable
	wire         seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_readdatavalid;                    // seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:av_readdatavalid -> seq_trk_mgr_inst_avl_translator:uav_readdatavalid
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // mmr_bridge_s0_translator:uav_waitrequest -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> mmr_bridge_s0_translator:uav_burstcount
	wire  [31:0] mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                             // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> mmr_bridge_s0_translator:uav_writedata
	wire  [19:0] mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                               // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> mmr_bridge_s0_translator:uav_address
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                                 // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> mmr_bridge_s0_translator:uav_write
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                  // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> mmr_bridge_s0_translator:uav_lock
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                                  // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> mmr_bridge_s0_translator:uav_read
	wire  [31:0] mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                              // mmr_bridge_s0_translator:uav_readdata -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // mmr_bridge_s0_translator:uav_readdatavalid -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mmr_bridge_s0_translator:uav_debugaccess
	wire   [3:0] mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> mmr_bridge_s0_translator:uav_byteenable
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [73:0] mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                           // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [73:0] mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // seq_scc_mgr_inst_avl_translator:uav_waitrequest -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:m0_burstcount -> seq_scc_mgr_inst_avl_translator:uav_burstcount
	wire  [31:0] seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_writedata;                // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:m0_writedata -> seq_scc_mgr_inst_avl_translator:uav_writedata
	wire  [19:0] seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_address;                  // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:m0_address -> seq_scc_mgr_inst_avl_translator:uav_address
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_write;                    // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:m0_write -> seq_scc_mgr_inst_avl_translator:uav_write
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_lock;                     // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:m0_lock -> seq_scc_mgr_inst_avl_translator:uav_lock
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_read;                     // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:m0_read -> seq_scc_mgr_inst_avl_translator:uav_read
	wire  [31:0] seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // seq_scc_mgr_inst_avl_translator:uav_readdata -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // seq_scc_mgr_inst_avl_translator:uav_readdatavalid -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> seq_scc_mgr_inst_avl_translator:uav_debugaccess
	wire   [3:0] seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:m0_byteenable -> seq_scc_mgr_inst_avl_translator:uav_byteenable
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rf_source_valid -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [73:0] seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_data;              // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rf_source_data -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [73:0] seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // hphy_bridge_s0_translator:uav_waitrequest -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> hphy_bridge_s0_translator:uav_burstcount
	wire  [31:0] hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                            // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> hphy_bridge_s0_translator:uav_writedata
	wire  [19:0] hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                              // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> hphy_bridge_s0_translator:uav_address
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                                // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> hphy_bridge_s0_translator:uav_write
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                 // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> hphy_bridge_s0_translator:uav_lock
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                                 // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> hphy_bridge_s0_translator:uav_read
	wire  [31:0] hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                             // hphy_bridge_s0_translator:uav_readdata -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // hphy_bridge_s0_translator:uav_readdatavalid -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hphy_bridge_s0_translator:uav_debugaccess
	wire   [3:0] hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> hphy_bridge_s0_translator:uav_byteenable
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [73:0] hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                          // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [73:0] hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                            // cpu_inst_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_valid;                                  // cpu_inst_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                          // cpu_inst_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [72:0] cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_data;                                   // cpu_inst_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_ready;                                  // addr_router:sink_ready -> cpu_inst_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire         seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_endofpacket;             // seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_valid;                   // seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_startofpacket;           // seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [72:0] seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_data;                    // seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_ready;                   // addr_router_001:sink_ready -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:cp_ready
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                 // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [72:0] mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                                  // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router:sink_ready -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                                // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [72:0] hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                                 // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_001:sink_ready -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_valid;                    // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [72:0] seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_data;                     // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_002:sink_ready -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_valid;                   // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [72:0] seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_data;                    // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_003:sink_ready -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                      // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                            // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                    // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [72:0] addr_router_src_data;                                                                             // addr_router:src_data -> limiter:cmd_sink_data
	wire   [3:0] addr_router_src_channel;                                                                          // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                            // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                      // limiter:rsp_src_endofpacket -> cpu_inst_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                            // limiter:rsp_src_valid -> cpu_inst_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                    // limiter:rsp_src_startofpacket -> cpu_inst_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [72:0] limiter_rsp_src_data;                                                                             // limiter:rsp_src_data -> cpu_inst_m0_translator_avalon_universal_master_0_agent:rp_data
	wire   [3:0] limiter_rsp_src_channel;                                                                          // limiter:rsp_src_channel -> cpu_inst_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                            // cpu_inst_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         cmd_xbar_demux_src0_endofpacket;                                                                  // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                        // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [72:0] cmd_xbar_demux_src0_data;                                                                         // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [3:0] cmd_xbar_demux_src0_channel;                                                                      // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                        // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                  // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                        // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [72:0] cmd_xbar_demux_src1_data;                                                                         // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [3:0] cmd_xbar_demux_src1_channel;                                                                      // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                        // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                  // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                        // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [72:0] cmd_xbar_demux_src2_data;                                                                         // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [3:0] cmd_xbar_demux_src2_channel;                                                                      // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                        // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_src3_endofpacket;                                                                  // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                        // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [72:0] cmd_xbar_demux_src3_data;                                                                         // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [3:0] cmd_xbar_demux_src3_channel;                                                                      // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire         cmd_xbar_demux_src3_ready;                                                                        // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                              // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                    // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                            // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [72:0] cmd_xbar_demux_001_src0_data;                                                                     // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [3:0] cmd_xbar_demux_001_src0_channel;                                                                  // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                    // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                              // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                    // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                            // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [72:0] cmd_xbar_demux_001_src1_data;                                                                     // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [3:0] cmd_xbar_demux_001_src1_channel;                                                                  // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                    // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                              // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                    // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                            // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [72:0] cmd_xbar_demux_001_src2_data;                                                                     // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [3:0] cmd_xbar_demux_001_src2_channel;                                                                  // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                    // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                              // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                    // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                            // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [72:0] cmd_xbar_demux_001_src3_data;                                                                     // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [3:0] cmd_xbar_demux_001_src3_channel;                                                                  // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire         cmd_xbar_demux_001_src3_ready;                                                                    // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                                  // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                        // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [72:0] rsp_xbar_demux_src0_data;                                                                         // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [3:0] rsp_xbar_demux_src0_channel;                                                                      // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                        // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                  // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                        // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [72:0] rsp_xbar_demux_src1_data;                                                                         // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [3:0] rsp_xbar_demux_src1_channel;                                                                      // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                        // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                              // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                    // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                            // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [72:0] rsp_xbar_demux_001_src0_data;                                                                     // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [3:0] rsp_xbar_demux_001_src0_channel;                                                                  // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                    // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                              // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                    // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                            // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [72:0] rsp_xbar_demux_001_src1_data;                                                                     // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [3:0] rsp_xbar_demux_001_src1_channel;                                                                  // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                    // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                              // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                    // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                            // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [72:0] rsp_xbar_demux_002_src0_data;                                                                     // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [3:0] rsp_xbar_demux_002_src0_channel;                                                                  // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                    // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                              // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                    // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                            // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [72:0] rsp_xbar_demux_002_src1_data;                                                                     // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [3:0] rsp_xbar_demux_002_src1_channel;                                                                  // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                    // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                              // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                    // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                            // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [72:0] rsp_xbar_demux_003_src0_data;                                                                     // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [3:0] rsp_xbar_demux_003_src0_channel;                                                                  // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                    // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_003_src1_endofpacket;                                                              // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src1_valid;                                                                    // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src1_startofpacket;                                                            // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [72:0] rsp_xbar_demux_003_src1_data;                                                                     // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [3:0] rsp_xbar_demux_003_src1_channel;                                                                  // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src1_ready;                                                                    // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire         limiter_cmd_src_endofpacket;                                                                      // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                    // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [72:0] limiter_cmd_src_data;                                                                             // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [3:0] limiter_cmd_src_channel;                                                                          // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                            // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                     // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                           // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                   // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [72:0] rsp_xbar_mux_src_data;                                                                            // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [3:0] rsp_xbar_mux_src_channel;                                                                         // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                           // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                  // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                        // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [72:0] addr_router_001_src_data;                                                                         // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [3:0] addr_router_001_src_channel;                                                                      // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                        // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                 // rsp_xbar_mux_001:src_endofpacket -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                       // rsp_xbar_mux_001:src_valid -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                               // rsp_xbar_mux_001:src_startofpacket -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [72:0] rsp_xbar_mux_001_src_data;                                                                        // rsp_xbar_mux_001:src_data -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:rp_data
	wire   [3:0] rsp_xbar_mux_001_src_channel;                                                                     // rsp_xbar_mux_001:src_channel -> seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                       // seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                     // cmd_xbar_mux:src_endofpacket -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                           // cmd_xbar_mux:src_valid -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                   // cmd_xbar_mux:src_startofpacket -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [72:0] cmd_xbar_mux_src_data;                                                                            // cmd_xbar_mux:src_data -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_mux_src_channel;                                                                         // cmd_xbar_mux:src_channel -> mmr_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                           // mmr_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                        // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                              // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                      // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [72:0] id_router_src_data;                                                                               // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [3:0] id_router_src_channel;                                                                            // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                              // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                 // cmd_xbar_mux_001:src_endofpacket -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                       // cmd_xbar_mux_001:src_valid -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                               // cmd_xbar_mux_001:src_startofpacket -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [72:0] cmd_xbar_mux_001_src_data;                                                                        // cmd_xbar_mux_001:src_data -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_mux_001_src_channel;                                                                     // cmd_xbar_mux_001:src_channel -> hphy_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                       // hphy_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                    // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                          // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                  // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [72:0] id_router_001_src_data;                                                                           // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [3:0] id_router_001_src_channel;                                                                        // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                          // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                 // cmd_xbar_mux_002:src_endofpacket -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                       // cmd_xbar_mux_002:src_valid -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                               // cmd_xbar_mux_002:src_startofpacket -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [72:0] cmd_xbar_mux_002_src_data;                                                                        // cmd_xbar_mux_002:src_data -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_mux_002_src_channel;                                                                     // cmd_xbar_mux_002:src_channel -> seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                       // seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                    // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                          // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                  // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [72:0] id_router_002_src_data;                                                                           // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [3:0] id_router_002_src_channel;                                                                        // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                          // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_mux_003_src_endofpacket;                                                                 // cmd_xbar_mux_003:src_endofpacket -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_003_src_valid;                                                                       // cmd_xbar_mux_003:src_valid -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_003_src_startofpacket;                                                               // cmd_xbar_mux_003:src_startofpacket -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [72:0] cmd_xbar_mux_003_src_data;                                                                        // cmd_xbar_mux_003:src_data -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:cp_data
	wire   [3:0] cmd_xbar_mux_003_src_channel;                                                                     // cmd_xbar_mux_003:src_channel -> seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_003_src_ready;                                                                       // seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire         id_router_003_src_endofpacket;                                                                    // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                          // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                  // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [72:0] id_router_003_src_data;                                                                           // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [3:0] id_router_003_src_channel;                                                                        // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                          // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire   [3:0] limiter_cmd_valid_data;                                                                           // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid







	assign scc_dqsb_ena = scc_dqs_ena;


	seq_altera_hhp_apb2avalon_bridge #(
		.DWIDTH           (32),
		.AWIDTH           (32),
		.BYTEENABLE_WIDTH (4)
	) apb2avalon_bridge_inst (
		.av_addr        (apb2avalon_bridge_inst_avalon_master_address),       // avalon_master.address
		.av_write       (apb2avalon_bridge_inst_avalon_master_write),         //              .write
		.av_read        (apb2avalon_bridge_inst_avalon_master_read),          //              .read
		.av_writedata   (apb2avalon_bridge_inst_avalon_master_writedata),     //              .writedata
		.av_readdata    (apb2avalon_bridge_inst_avalon_master_readdata),      //              .readdata
		.av_rdata_valid (apb2avalon_bridge_inst_avalon_master_readdatavalid), //              .readdatavalid
		.av_byteenable  (apb2avalon_bridge_inst_avalon_master_byteenable),    //              .byteenable
		.av_waitrequest (apb2avalon_bridge_inst_avalon_master_waitrequest),   //              .waitrequest
		.prdata         (prdata),                                             //     apb_slave.prdata
		.pready         (pready),                                             //              .pready
		.pslverr        (pslverr),                                            //              .pslverr
		.pwdata         (pwdata),                                             //              .pwdata
		.pwrite         (pwrite),                                             //              .pwrite
		.penable        (penable),                                            //              .penable
		.psel           (psel),                                               //              .psel
		.paddr          (paddr),                                              //              .paddr
		.clk_p           (apb_clk),                                            //          pclk.clk
		.sp_reset_n     (apb_reset_n),                    		      //    sp_reset_n.reset_n
		.debug_hphy_reg (debug_hphy_reg_apb2avl), 
		.debug_hphy_comb(debug_hphy_comb_apb2avl)

	);

	seq_altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (20),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) cpu_inst (
		.m0_clk           (avl_clk),                                                  //   m0_clk.clk
		.m0_reset_n       (avl_reset_n),                       // m0_reset.reset
		.s0_clk           (apb_clk),                                                  //   s0_clk.clk
		.s0_reset_n       (apb_reset_n),                           // s0_reset.reset
		.s0_waitrequest   (cpu_inst_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (cpu_inst_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (cpu_inst_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (cpu_inst_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (cpu_inst_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (cpu_inst_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (cpu_inst_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (cpu_inst_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (cpu_inst_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (cpu_inst_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (cpu_inst_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (cpu_inst_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (cpu_inst_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (cpu_inst_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (cpu_inst_m0_writedata),                                    //         .writedata
		.m0_address       (cpu_inst_m0_address),                                      //         .address
		.m0_write         (cpu_inst_m0_write),                                        //         .write
		.m0_read          (cpu_inst_m0_read),                                         //         .read
		.m0_byteenable    (cpu_inst_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (cpu_inst_m0_debugaccess),                                  //         .debugaccess
		.debug_hphy_reg   (debug_hphy_reg_clk_crossing), 
		.debug_hphy_comb  (debug_hphy_comb_clk_crossing)
		
	);

	seq_hhp_decompress_avl_mm_bridge #(
		.DATA_WIDTH    (32),
		.SYMBOL_WIDTH  (8),
		.ADDRESS_WIDTH (32)
	) seq_hhp_decompress_bridge (
		.clk              (apb_clk),                                                             //   clk.clk
		.reset_n          (apb_reset_n),                                     // reset.reset_n
		.s0_address       (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_address),     //    s0.address
		.s0_read          (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_read),        //      .read
		.s0_readdata      (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_readdata),    //      .readdata
		.s0_write         (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_write),       //      .write
		.s0_writedata     (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_writedata),   //      .writedata
		.s0_waitrequest   (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_waitrequest), //      .waitrequest
		.m0_address       (seq_hhp_decompress_bridge_m0_address),                                    //    m0.address
		.m0_read          (seq_hhp_decompress_bridge_m0_read),                                       //      .read
		.m0_readdata      (seq_hhp_decompress_bridge_m0_readdata),                                   //      .readdata
		.m0_write         (seq_hhp_decompress_bridge_m0_write),                                      //      .write
		.m0_writedata     (seq_hhp_decompress_bridge_m0_writedata),                                  //      .writedata
		.m0_waitrequest   (seq_hhp_decompress_bridge_m0_waitrequest),                                //      .waitrequest
		.s0_byteenable    (4'b1111),                                                             // (terminated)
		.s0_readdatavalid (),                                                                    // (terminated)
		.m0_byteenable    (),                                                                    // (terminated)
		.m0_readdatavalid (1'b0),                                                                 // (terminated)
		.debug_hphy_comb  (debug_hphy_comb_decompress)
		
	);

	seq_altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (8),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mmr_bridge (
		.clk              (avl_clk),                                                    //   clk.clk
		.reset_n          (avl_reset_n),                         // reset.reset
		.s0_waitrequest   (mmr_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mmr_bridge_s0_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.s0_readdatavalid (mmr_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mmr_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.s0_writedata     (mmr_bridge_s0_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.s0_address       (mmr_bridge_s0_translator_avalon_anti_slave_0_address),       //      .address
		.s0_write         (mmr_bridge_s0_translator_avalon_anti_slave_0_write),         //      .write
		.s0_read          (mmr_bridge_s0_translator_avalon_anti_slave_0_read),          //      .read
		.s0_byteenable    (mmr_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.s0_debugaccess   (mmr_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mmr_avl_waitrequest),                                        //    m0.waitrequest
		.m0_readdata      (mmr_avl_readdata),                                           //      .readdata
		.m0_readdatavalid (mmr_avl_readdatavalid),                                      //      .readdatavalid
		.m0_burstcount    (mmr_avl_burstcount),                                         //      .burstcount
		.m0_writedata     (mmr_avl_writedata),                                          //      .writedata
		.m0_address       (mmr_avl_address),                                            //      .address
		.m0_write         (mmr_avl_write),                                              //      .write
		.m0_read          (mmr_avl_read),                                               //      .read
//		.m0_byteenable    (mmr_avl_be),                                                 //      .byteenable
		.m0_debugaccess   (mmr_avl_debugaccess)                                         //      .debugaccess
	);

	seq_scc_mgr #(
		.AVL_DATA_WIDTH         (32),
		.AVL_ADDR_WIDTH         (13),
		.MEM_IF_READ_DQS_WIDTH  (5),
		.MEM_IF_WRITE_DQS_WIDTH (5),
		.MEM_IF_DQ_WIDTH        (40),
		.MEM_IF_DM_WIDTH        (5),
		.DLL_DELAY_CHAIN_LENGTH (8),
		.HHP_HPS                (1),
		.DQS_TRK_ENABLED        (1),
		.DUAL_WRITE_CLOCK       (0)
	) seq_scc_mgr_inst (
		.avl_clk                 (avl_clk),                                                               //          avl_clk.clk
		.avl_reset_n             (avl_reset_n),                                   //        avl_reset.reset_n
		.avl_address             (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_address),     //              avl.address
		.avl_write               (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_write),       //                 .write
		.avl_writedata           (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_writedata),   //                 .writedata
		.avl_read                (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_read),        //                 .read
		.avl_readdata            (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_readdata),    //                 .readdata
		.avl_waitrequest         (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_waitrequest), //                 .waitrequest
		.scc_clk                 (avl_clk),                                                               //          scc_clk.clk
		.scc_clk_out             (scc_clk_out),
		.scc_reset_n             (avl_reset_n),
		.scc_data                (scc_data),                                                              //              scc.scc_data
		.scc_dqs_ena             (scc_dqs_ena),                                                           //                 .scc_dqs_ena
		.scc_dqs_io_ena          (scc_dqs_io_ena),                                                        //                 .scc_dqs_io_ena
		.scc_dq_ena              (scc_dq_ena),                                                            //                 .scc_dq_ena
		.scc_dm_ena              (scc_dm_ena),                                                            //                 .scc_dm_ena
		.scc_upd                 (scc_upd),                                                               //                 .scc_upd
		.capture_strobe_tracking (capture_strobe_tracking),                                               //                 .capture_strobe_tracking
		.afi_init_req            (afi_init_req),                                                          // afi_init_cal_req.afi_init_req
		.afi_cal_req             (afi_cal_req),                                                            //                 .afi_cal_req
		.debug_hphy_reg		 (debug_hphy_reg_scc), 
		.debug_hphy_comb	 (debug_hphy_comb_scc)
	);

	seq_reg_file #(
		.AVL_DATA_WIDTH    (32),
		.AVL_ADDR_WIDTH    (13),
		.AVL_NUM_SYMBOLS   (4),
		.AVL_SYMBOL_WIDTH  (8),
		.REGISTER_RDATA    (0),
		.NUM_REGFILE_WORDS (16)
	) seq_reg_file_inst (
		.avl_clk         (avl_clk),                                                                //   avl_clk.clk
		.avl_reset_n     (avl_reset_n),                                    // avl_reset.reset_n
		.avl_address     (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_address),     //       avl.address
		.avl_write       (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_write),       //          .write
		.avl_writedata   (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_writedata),   //          .writedata
		.avl_read        (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_read),        //          .read
		.avl_readdata    (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_readdata),    //          .readdata
		.avl_waitrequest (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_waitrequest), //          .waitrequest
		.avl_be          (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_byteenable),  //          .byteenable
		.debug_hphy_reg  (debug_hphy_reg_reg), 
		.debug_hphy_comb (debug_hphy_comb_reg)

	);

	seq_altera_mem_if_simple_avalon_mm_bridge #(
		.DATA_WIDTH                (32),
		.SYMBOL_WIDTH              (8),
		.ADDRESS_WIDTH             (16)
	) hphy_bridge (
		.clk              (avl_clk),                                                   //   clk.clk
		.reset_n          (avl_reset_n),                       // reset.reset_n
		.s0_address       (hphy_bridge_s0_translator_avalon_anti_slave_0_address),     //    s0.address
		.s0_read          (hphy_bridge_s0_translator_avalon_anti_slave_0_read),        //      .read
		.s0_readdata      (hphy_bridge_s0_translator_avalon_anti_slave_0_readdata),    //      .readdata
		.s0_write         (hphy_bridge_s0_translator_avalon_anti_slave_0_write),       //      .write
		.s0_writedata     (hphy_bridge_s0_translator_avalon_anti_slave_0_writedata),   //      .writedata
		.s0_waitrequest   (hphy_bridge_s0_translator_avalon_anti_slave_0_waitrequest), //      .waitrequest
		.m0_address       (avl_address),                                               //    m0.address
		.m0_read          (avl_read),                                                  //      .read
		.m0_readdata      (avl_readdata),                                              //      .readdata
		.m0_write         (avl_write),                                                 //      .write
		.m0_writedata     (avl_writedata),                                             //      .writedata
		.m0_waitrequest   (avl_waitrequest),                                           //      .waitrequest
		.s0_byteenable    (4'b1111),                                                   // (terminated)
		.s0_readdatavalid (),                                                          // (terminated)
		.m0_byteenable    (),                                                          // (terminated)
		.m0_readdatavalid (1'b0)                                                       // (terminated)
	);

	seq_trk_mgr #(
		.MEM_CHIP_SELECT_WIDTH  (2),
		.AVL_DATA_WIDTH         (32),
		.AVL_MTR_ADDR_WIDTH     (20),
		.MEM_DQS_WIDTH          (5),
		.PHASE_WIDTH            (3),
		.READ_VALID_FIFO_SIZE   (16),
		.MUX_SEL_SEQUENCER_VAL  (3),
		.MUX_SEL_CONTROLLER_VAL (2),
		.PHY_MGR_BASE           (557056),
		.RW_MGR_BASE            (589824),
		.SCC_MGR_BASE           (65536),
		.REG_FILE_BASE          (98304)
	) seq_trk_mgr_inst (
		.avl_clk              (avl_clk),                                //   avl_clk.clk
		.avl_reset_n          (avl_reset_n),    // avl_reset.reset_n
		.avl_address          (seq_trk_mgr_inst_avl_address),     //       avl.address
		.avl_write            (seq_trk_mgr_inst_avl_write),       //          .write
		.avl_writedata        (seq_trk_mgr_inst_avl_writedata),   //          .writedata
		.avl_read             (seq_trk_mgr_inst_avl_read),        //          .read
		.avl_readdata         (seq_trk_mgr_inst_avl_readdata),    //          .readdata
		.avl_waitrequest      (seq_trk_mgr_inst_avl_waitrequest), //          .waitrequest
		.afi_seq_busy         (afi_seq_busy),                           //       afi.afi_seq_busy
		.afi_ctl_long_idle    (afi_ctl_long_idle),                      //          .afi_ctl_long_idle
		.afi_ctl_refresh_done (afi_ctl_refresh_done),                    //          .afi_ctl_refresh_done
		.debug_hphy_reg	      (debug_hphy_reg_trck), 
		.debug_hphy_comb      (debug_hphy_comb_trck)
	);

	seq_altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (1),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) apb2avalon_bridge_inst_avalon_master_translator (
		.clk                   (apb_clk),                                                                                 //                       clk.clk
		.reset_n               (apb_reset_n),                                                          //                     reset.reset
		.uav_address           (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (apb2avalon_bridge_inst_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (apb2avalon_bridge_inst_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (apb2avalon_bridge_inst_avalon_master_byteenable),                                         //                          .byteenable
		.av_read               (apb2avalon_bridge_inst_avalon_master_read),                                               //                          .read
		.av_readdata           (apb2avalon_bridge_inst_avalon_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (apb2avalon_bridge_inst_avalon_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (apb2avalon_bridge_inst_avalon_master_write),                                              //                          .write
		.av_writedata          (apb2avalon_bridge_inst_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                                    //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                    //               (terminated)
		.av_begintransfer      (1'b0),                                                                                    //               (terminated)
		.av_chipselect         (1'b0),                                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                                    //               (terminated)
		.av_debugaccess        (1'b0),                                                                                    //               (terminated)
		.uav_clken             (),                                                                                        //               (terminated)
		.av_clken              (1'b1)                                                                                     //               (terminated)
	);

	seq_altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (32),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) seq_hhp_decompress_bridge_s0_translator (
		.clk                   (apb_clk),                                                                                 //                      clk.clk
		.reset_n               (apb_reset_n),                                                          //                    reset.reset
		.uav_address           (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read              (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write             (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest       (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata          (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata         (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock              (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess       (apb2avalon_bridge_inst_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address            (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_address),                         //      avalon_anti_slave_0.address
		.av_write              (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_write),                           //                         .write
		.av_read               (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_read),                            //                         .read
		.av_readdata           (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_readdata),                        //                         .readdata
		.av_writedata          (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_writedata),                       //                         .writedata
		.av_waitrequest        (seq_hhp_decompress_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                     //                         .waitrequest
		.av_begintransfer      (),                                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                                        //              (terminated)
		.av_burstcount         (),                                                                                        //              (terminated)
		.av_byteenable         (),                                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                        //              (terminated)
		.av_lock               (),                                                                                        //              (terminated)
		.av_chipselect         (),                                                                                        //              (terminated)
		.av_clken              (),                                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                                    //              (terminated)
		.av_debugaccess        (),                                                                                        //              (terminated)
		.av_outputenable       ()                                                                                         //              (terminated)
	);

	seq_altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) seq_hhp_decompress_bridge_m0_translator (
		.clk                   (apb_clk),                                                                     //                       clk.clk
		.reset_n               (apb_reset_n),                                              //                     reset.reset
		.uav_address           (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (seq_hhp_decompress_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (seq_hhp_decompress_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_read               (seq_hhp_decompress_bridge_m0_read),                                               //                          .read
		.av_readdata           (seq_hhp_decompress_bridge_m0_readdata),                                           //                          .readdata
		.av_write              (seq_hhp_decompress_bridge_m0_write),                                              //                          .write
		.av_writedata          (seq_hhp_decompress_bridge_m0_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_readdatavalid      (),                                                                            //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	seq_altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (20),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_inst_s0_translator (
		.clk                   (apb_clk),                                                                     //                      clk.clk
		.reset_n               (apb_reset_n),                                              //                    reset.reset
		.uav_address           (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read              (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write             (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest       (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata          (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata         (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock              (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess       (seq_hhp_decompress_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address            (cpu_inst_s0_translator_avalon_anti_slave_0_address),                          //      avalon_anti_slave_0.address
		.av_write              (cpu_inst_s0_translator_avalon_anti_slave_0_write),                            //                         .write
		.av_read               (cpu_inst_s0_translator_avalon_anti_slave_0_read),                             //                         .read
		.av_readdata           (cpu_inst_s0_translator_avalon_anti_slave_0_readdata),                         //                         .readdata
		.av_writedata          (cpu_inst_s0_translator_avalon_anti_slave_0_writedata),                        //                         .writedata
		.av_burstcount         (cpu_inst_s0_translator_avalon_anti_slave_0_burstcount),                       //                         .burstcount
		.av_byteenable         (cpu_inst_s0_translator_avalon_anti_slave_0_byteenable),                       //                         .byteenable
		.av_readdatavalid      (cpu_inst_s0_translator_avalon_anti_slave_0_readdatavalid),                    //                         .readdatavalid
		.av_waitrequest        (cpu_inst_s0_translator_avalon_anti_slave_0_waitrequest),                      //                         .waitrequest
		.av_debugaccess        (cpu_inst_s0_translator_avalon_anti_slave_0_debugaccess),                      //                         .debugaccess
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_chipselect         (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	seq_altera_merlin_master_translator #(
		.AV_ADDRESS_W                (20),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (20),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_inst_m0_translator (
		.clk                   (avl_clk),                                                        //                       clk.clk
		.reset_n               (avl_reset_n),                             //                     reset.reset
		.uav_address           (cpu_inst_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_inst_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_inst_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_inst_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_inst_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_inst_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_inst_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_inst_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_inst_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_inst_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_inst_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_inst_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_inst_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (cpu_inst_m0_burstcount),                                         //                          .burstcount
		.av_byteenable         (cpu_inst_m0_byteenable),                                         //                          .byteenable
		.av_read               (cpu_inst_m0_read),                                               //                          .read
		.av_readdata           (cpu_inst_m0_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_inst_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (cpu_inst_m0_write),                                              //                          .write
		.av_writedata          (cpu_inst_m0_writedata),                                          //                          .writedata
		.av_debugaccess        (cpu_inst_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer (1'b0),                                                           //               (terminated)
		.av_begintransfer      (1'b0),                                                           //               (terminated)
		.av_chipselect         (1'b0),                                                           //               (terminated)
		.av_lock               (1'b0),                                                           //               (terminated)
		.uav_clken             (),                                                               //               (terminated)
		.av_clken              (1'b1)                                                            //               (terminated)
	);

	seq_altera_merlin_master_translator #(
		.AV_ADDRESS_W                (20),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (20),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) seq_trk_mgr_inst_avl_translator (
		.clk                   (avl_clk),                                                                       //                       clk.clk
		.reset_n               (avl_reset_n),                                            //                     reset.reset
		.uav_address           (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (seq_trk_mgr_inst_avl_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (seq_trk_mgr_inst_avl_waitrequest),                                        //                          .waitrequest
		.av_read               (seq_trk_mgr_inst_avl_read),                                               //                          .read
		.av_readdata           (seq_trk_mgr_inst_avl_readdata),                                           //                          .readdata
		.av_write              (seq_trk_mgr_inst_avl_write),                                              //                          .write
		.av_writedata          (seq_trk_mgr_inst_avl_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                          //               (terminated)
		.av_byteenable         (4'b1111),                                                                       //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                          //               (terminated)
		.av_begintransfer      (1'b0),                                                                          //               (terminated)
		.av_chipselect         (1'b0),                                                                          //               (terminated)
		.av_readdatavalid      (),                                                                              //               (terminated)
		.av_lock               (1'b0),                                                                          //               (terminated)
		.av_debugaccess        (1'b0),                                                                          //               (terminated)
		.uav_clken             (),                                                                              //               (terminated)
		.av_clken              (1'b1)                                                                           //               (terminated)
	);

	seq_altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mmr_bridge_s0_translator (
		.clk                   (avl_clk),                                                                  //                      clk.clk
		.reset_n               (avl_reset_n),                                       //                    reset.reset
		.uav_address           (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (mmr_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (mmr_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (mmr_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (mmr_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (mmr_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (mmr_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (mmr_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (mmr_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (mmr_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess        (mmr_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_chipselect         (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	seq_altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (16),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hphy_bridge_s0_translator (
		.clk                   (avl_clk),                                                                   //                      clk.clk
		.reset_n               (avl_reset_n),                                        //                    reset.reset
		.uav_address           (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (hphy_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (hphy_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (hphy_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (hphy_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (hphy_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (hphy_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_byteenable         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_chipselect         (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	seq_altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) seq_scc_mgr_inst_avl_translator (
		.clk                   (avl_clk),                                                                               //                      clk.clk
		.reset_n               (avl_reset_n),                                                    //                    reset.reset
		.uav_address           (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (seq_scc_mgr_inst_avl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                      //              (terminated)
		.av_byteenable         (),                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                      //              (terminated)
		.av_lock               (),                                                                                      //              (terminated)
		.av_chipselect         (),                                                                                      //              (terminated)
		.av_clken              (),                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                       //              (terminated)
	);

	seq_altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (20),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) seq_reg_file_inst_avl_translator (
		.clk                   (avl_clk),                                                                                //                      clk.clk
		.reset_n               (avl_reset_n),                                                     //                    reset.reset
		.uav_address           (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (seq_reg_file_inst_avl_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_chipselect         (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	seq_altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (67),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (72),
		.PKT_PROTECTION_L          (72),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (73),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent (
		.clk                     (avl_clk),                                                                                          //             clk.clk
		.reset_n                 (avl_reset_n),                                                               //       clk_reset.reset
		.m0_address              (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                                     //                .channel
		.rf_sink_ready           (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	seq_altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (74),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (avl_clk),                                                                                          //       clk.clk
		.reset_n           (avl_reset_n),                                                               // clk_reset.reset
		.in_data           (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	seq_altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (72),
		.PKT_PROTECTION_L          (72),
		.PKT_BEGIN_BURST           (67),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.ST_DATA_W                 (73),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7)
	) cpu_inst_m0_translator_avalon_universal_master_0_agent (
		.clk              (avl_clk),                                                                 //       clk.clk
		.reset_n          (~avl_reset_n),                                      // clk_reset.reset
		.av_address       (cpu_inst_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_inst_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_inst_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_inst_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_inst_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_inst_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_inst_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_inst_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_inst_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_inst_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_inst_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                   //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                    //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                 //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                             //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                    //          .ready
	);

	seq_altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (72),
		.PKT_PROTECTION_L          (72),
		.PKT_BEGIN_BURST           (67),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.ST_DATA_W                 (73),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7)
	) seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent (
		.clk              (avl_clk),                                                                                //       clk.clk
		.reset_n          (avl_reset_n),                                                     // clk_reset.reset
		.av_address       (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                             //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                              //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                           //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                                       //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                              //          .ready
	);

	seq_altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (67),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (72),
		.PKT_PROTECTION_L          (72),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (73),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) mmr_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (avl_clk),                                                                            //             clk.clk
		.reset_n                 (avl_reset_n),                                                 //       clk_reset.reset
		.m0_address              (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                           //                .channel
		.rf_sink_ready           (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	seq_altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (74),
		.FIFO_DEPTH          (5),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (avl_clk),                                                                            //       clk.clk
		.reset_n           (avl_reset_n),                                                 // clk_reset.reset
		.in_data           (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	seq_altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (67),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (72),
		.PKT_PROTECTION_L          (72),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (73),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent (
		.clk                     (avl_clk),                                                                                         //             clk.clk
		.reset_n                 (avl_reset_n),                                                              //       clk_reset.reset
		.m0_address              (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                                    //                .channel
		.rf_sink_ready           (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	seq_altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (74),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (avl_clk),                                                                                         //       clk.clk
		.reset_n           (avl_reset_n),                                                              // clk_reset.reset
		.in_data           (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	seq_altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (67),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (55),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (56),
		.PKT_TRANS_POSTED          (57),
		.PKT_TRANS_WRITE           (58),
		.PKT_TRANS_READ            (59),
		.PKT_TRANS_LOCK            (60),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (68),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_PROTECTION_H          (72),
		.PKT_PROTECTION_L          (72),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (73),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) hphy_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (avl_clk),                                                                             //             clk.clk
		.reset_n                 (avl_reset_n),                                                  //       clk_reset.reset
		.m0_address              (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                        //                .channel
		.rf_sink_ready           (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	seq_altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (74),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (avl_clk),                                                                             //       clk.clk
		.reset_n           (avl_reset_n),                                                  // clk_reset.reset
		.in_data           (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	seq_addr_router addr_router (
		.sink_ready         (cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_inst_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (avl_clk),                                                                 //       clk.clk
		.reset_n            (avl_reset_n),                                      // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_src_valid),                                                   //          .valid
		.src_data           (addr_router_src_data),                                                    //          .data
		.src_channel        (addr_router_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                              //          .endofpacket
	);

	seq_addr_router_001 addr_router_001 (
		.sink_ready         (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (seq_trk_mgr_inst_avl_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (avl_clk),                                                                                //       clk.clk
		.reset_n            (avl_reset_n),                                                     // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                              //          .valid
		.src_data           (addr_router_001_src_data),                                                               //          .data
		.src_channel        (addr_router_001_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                         //          .endofpacket
	);

	seq_id_router id_router (
		.sink_ready         (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mmr_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (avl_clk),                                                                  //       clk.clk
		.reset_n            (avl_reset_n),                                       // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                      //       src.ready
		.src_valid          (id_router_src_valid),                                                      //          .valid
		.src_data           (id_router_src_data),                                                       //          .data
		.src_channel        (id_router_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                 //          .endofpacket
	);

	seq_id_router id_router_001 (
		.sink_ready         (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hphy_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (avl_clk),                                                                   //       clk.clk
		.reset_n            (avl_reset_n),                                        // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                   //       src.ready
		.src_valid          (id_router_001_src_valid),                                                   //          .valid
		.src_data           (id_router_001_src_data),                                                    //          .data
		.src_channel        (id_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                              //          .endofpacket
	);

	seq_id_router id_router_002 (
		.sink_ready         (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (seq_scc_mgr_inst_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (avl_clk),                                                                               //       clk.clk
		.reset_n            (avl_reset_n),                                                    // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                               //       src.ready
		.src_valid          (id_router_002_src_valid),                                                               //          .valid
		.src_data           (id_router_002_src_data),                                                                //          .data
		.src_channel        (id_router_002_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                          //          .endofpacket
	);

	seq_id_router id_router_003 (
		.sink_ready         (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (seq_reg_file_inst_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (avl_clk),                                                                                //       clk.clk
		.reset_n            (avl_reset_n),                                                     // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                //          .valid
		.src_data           (id_router_003_src_data),                                                                 //          .data
		.src_channel        (id_router_003_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                           //          .endofpacket
	);

	seq_altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (70),
		.PKT_TRANS_POSTED          (57),
		.MAX_OUTSTANDING_RESPONSES (4),
		.PIPELINED                 (0),
		.ST_DATA_W                 (73),
		.ST_CHANNEL_W              (4),
		.VALID_WIDTH               (4),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (61),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (avl_clk),                            //       clk.clk
		.reset_n                (avl_reset_n), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),              //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),              //          .valid
		.cmd_sink_data          (addr_router_src_data),               //          .data
		.cmd_sink_channel       (addr_router_src_channel),            //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),             //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),             //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),           //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),              //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket),     //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),       //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	seq_cmd_xbar_demux cmd_xbar_demux (
		.clk                (avl_clk),                            //        clk.clk
		.reset_n            (avl_reset_n), //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),            //           .channel
		.sink_data          (limiter_cmd_src_data),               //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),    //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),          //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),          //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),           //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),        //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),    //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),          //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),          //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),           //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),        //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)     //           .endofpacket
	);

	seq_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (avl_clk),                               //       clk.clk
		.reset_n            (avl_reset_n),    // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	seq_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (avl_clk),                               //       clk.clk
		.reset_n             (avl_reset_n),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	seq_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (avl_clk),                               //       clk.clk
		.reset_n             (avl_reset_n),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	seq_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (avl_clk),                               //       clk.clk
		.reset_n             (avl_reset_n),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	seq_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (avl_clk),                               //       clk.clk
		.reset_n             (avl_reset_n),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	seq_rsp_xbar_demux rsp_xbar_demux (
		.clk                (avl_clk),                            //       clk.clk
		.reset_n            (avl_reset_n), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	seq_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (avl_clk),                               //       clk.clk
		.reset_n            (avl_reset_n),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	seq_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (avl_clk),                               //       clk.clk
		.reset_n            (avl_reset_n),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	seq_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (avl_clk),                               //       clk.clk
		.reset_n            (avl_reset_n),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	seq_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (avl_clk),                               //       clk.clk
		.reset_n             (avl_reset_n),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	seq_rsp_xbar_mux rsp_xbar_mux_001 (
		.clk                 (avl_clk),                               //       clk.clk
		.reset_n             (avl_reset_n),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	//debug signals
	assign debug_hphy_reg  = {debug_hphy_reg_scc,debug_hphy_reg_reg,debug_hphy_reg_trck,debug_hphy_reg_apb2avl,debug_hphy_reg_clk_crossing};
	assign debug_hphy_comb = {debug_hphy_comb_scc,debug_hphy_comb_reg,debug_hphy_comb_trck,debug_hphy_comb_apb2avl,debug_hphy_comb_decompress,debug_hphy_comb_clk_crossing};

endmodule
